##
## LEF for PtnCells ;
## created by Innovus v20.11-s130_1 on Fri Jan 17 11:01:24 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BATCHARGERcore
  CLASS BLOCK ;
  SIZE 850.000000 BY 320.000000 ;
  FOREIGN BATCHARGERcore 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN iforcedbat
    DIRECTION OUTPUT ;
    USE ANALOG ;
    PORT
      LAYER metal4 ;
        RECT 40.100000 0.000000 40.300000 0.520000 ;
    END
  END iforcedbat
  PIN vsensbat
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER metal4 ;
        RECT 200.100000 0.000000 200.300000 0.520000 ;
    END
  END vsensbat
  PIN vin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 849.360000 319.320000 850.000000 319.480000 ;
    END
  END vin
  PIN vbattemp
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER metal4 ;
        RECT 120.100000 0.000000 120.300000 0.520000 ;
    END
  END vbattemp
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 849.360000 212.920000 850.000000 213.080000 ;
    END
  END en
  PIN sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 849.360000 159.720000 850.000000 159.880000 ;
    END
  END sel[3]
  PIN sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 849.360000 106.520000 850.000000 106.680000 ;
    END
  END sel[2]
  PIN sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 849.360000 53.320000 850.000000 53.480000 ;
    END
  END sel[1]
  PIN sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 849.360000 0.120000 850.000000 0.280000 ;
    END
  END sel[0]
  PIN pgnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 849.360000 266.120000 850.000000 266.280000 ;
    END
  END pgnd
  PIN dvdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal3 ;
        RECT 424.500000 319.480000 424.700000 320.000000 ;
    END
  END dvdd
  PIN dgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal3 ;
        RECT 20.100000 319.480000 20.300000 320.000000 ;
    END
  END dgnd
  OBS
    LAYER metal1 ;
      RECT 0.000000 319.640000 850.000000 320.000000 ;
      RECT 0.000000 319.160000 849.170000 319.640000 ;
      RECT 0.000000 266.440000 850.000000 319.160000 ;
      RECT 0.000000 265.960000 849.170000 266.440000 ;
      RECT 0.000000 213.240000 850.000000 265.960000 ;
      RECT 0.000000 212.760000 849.170000 213.240000 ;
      RECT 0.000000 160.040000 850.000000 212.760000 ;
      RECT 0.000000 159.560000 849.170000 160.040000 ;
      RECT 0.000000 106.840000 850.000000 159.560000 ;
      RECT 0.000000 106.360000 849.170000 106.840000 ;
      RECT 0.000000 53.640000 850.000000 106.360000 ;
      RECT 0.000000 53.160000 849.170000 53.640000 ;
      RECT 0.000000 0.440000 850.000000 53.160000 ;
      RECT 0.000000 0.000000 849.170000 0.440000 ;
    LAYER metal2 ;
      RECT 0.000000 0.000000 850.000000 320.000000 ;
    LAYER metal3 ;
      RECT 424.900000 319.280000 850.000000 320.000000 ;
      RECT 20.500000 319.280000 424.300000 320.000000 ;
      RECT 0.000000 319.280000 19.900000 320.000000 ;
      RECT 0.000000 0.000000 850.000000 319.280000 ;
    LAYER metal4 ;
      RECT 0.000000 0.720000 850.000000 320.000000 ;
      RECT 200.500000 0.000000 850.000000 0.720000 ;
      RECT 120.500000 0.000000 199.900000 0.720000 ;
      RECT 40.500000 0.000000 119.900000 0.720000 ;
      RECT 0.000000 0.000000 39.900000 0.720000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 850.000000 320.000000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 850.000000 320.000000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 850.000000 320.000000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 850.000000 320.000000 ;
  END
END BATCHARGERcore

END LIBRARY
